-- megafunction wizard: %ALTIOBUF%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altiobuf_in 

-- ============================================================
-- File Name: ibuf.vhd
-- Megafunction Name(s):
-- 			altiobuf_in
--
-- Simulation Library Files(s):
-- 			cyclonev
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 16.1.0 Build 196 10/24/2016 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2016  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Intel and sold by Intel or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


--altiobuf_in CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" ENABLE_BUS_HOLD="FALSE" NUMBER_OF_CHANNELS=10 USE_DIFFERENTIAL_MODE="FALSE" USE_DYNAMIC_TERMINATION_CONTROL="TRUE" datain dataout
--VERSION_BEGIN 16.1 cbx_altiobuf_in 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_stratixiii 2016:10:24:15:04:16:SJ cbx_stratixv 2016:10:24:15:04:16:SJ  VERSION_END

 LIBRARY cyclonev;
 USE cyclonev.all;

--synthesis_resources = cyclonev_io_ibuf 10 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ibuf_iobuf_in_40i IS 
	 PORT 
	 ( 
		 datain	:	IN  STD_LOGIC_VECTOR (9 DOWNTO 0);
		 dataout	:	OUT  STD_LOGIC_VECTOR (9 DOWNTO 0)
	 ); 
 END ibuf_iobuf_in_40i;

 ARCHITECTURE RTL OF ibuf_iobuf_in_40i IS

	 SIGNAL  wire_ibufa_i	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_ibufa_o	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 COMPONENT  cyclonev_io_ibuf
	 GENERIC 
	 (
		bus_hold	:	STRING := "false";
		differential_mode	:	STRING := "false";
		simulate_z_as	:	STRING := "z";
		lpm_type	:	STRING := "cyclonev_io_ibuf"
	 );
	 PORT
	 ( 
		dynamicterminationcontrol	:	IN STD_LOGIC := '0';
		i	:	IN STD_LOGIC := '0';
		ibar	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	dataout <= wire_ibufa_o;
	wire_ibufa_i <= datain;
	loop0 : FOR i IN 0 TO 9 GENERATE 
	  ibufa :  cyclonev_io_ibuf
	  GENERIC MAP (
		bus_hold => "false",
		differential_mode => "false"
	  )
	  PORT MAP ( 
		i => wire_ibufa_i(i),
		o => wire_ibufa_o(i)
	  );
	END GENERATE loop0;

 END RTL; --ibuf_iobuf_in_40i
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ibuf IS
	PORT
	(
		datain		: IN STD_LOGIC_VECTOR (9 DOWNTO 0);
		dataout		: OUT STD_LOGIC_VECTOR (9 DOWNTO 0)
	);
END ibuf;


ARCHITECTURE RTL OF ibuf IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (9 DOWNTO 0);



	COMPONENT ibuf_iobuf_in_40i
	PORT (
			datain	: IN STD_LOGIC_VECTOR (9 DOWNTO 0);
			dataout	: OUT STD_LOGIC_VECTOR (9 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	dataout    <= sub_wire0(9 DOWNTO 0);

	ibuf_iobuf_in_40i_component : ibuf_iobuf_in_40i
	PORT MAP (
		datain => datain,
		dataout => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: enable_bus_hold STRING "FALSE"
-- Retrieval info: CONSTANT: number_of_channels NUMERIC "10"
-- Retrieval info: CONSTANT: use_differential_mode STRING "FALSE"
-- Retrieval info: CONSTANT: use_dynamic_termination_control STRING "TRUE"
-- Retrieval info: USED_PORT: datain 0 0 10 0 INPUT NODEFVAL "datain[9..0]"
-- Retrieval info: USED_PORT: dataout 0 0 10 0 OUTPUT NODEFVAL "dataout[9..0]"
-- Retrieval info: CONNECT: @datain 0 0 10 0 datain 0 0 10 0
-- Retrieval info: CONNECT: dataout 0 0 10 0 @dataout 0 0 10 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL ibuf.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ibuf.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ibuf.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ibuf.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ibuf_inst.vhd TRUE
-- Retrieval info: LIB_FILE: cyclonev
