library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package ov5640_controller_pkg is

	constant ov5640_init_wr_seq_len : integer := 211;
	type ov5640_init_wr_seq_t is array(0 to ov5640_init_wr_seq_len-1) of std_logic_vector(23 downto 0);
	
	constant ov5640_init_wr_seq : ov5640_init_wr_seq_t := (
	0   => x"3008" & x"82",
	1   => x"3008" & x"42",
	2   => x"3103" & x"03",
	3   => x"3017" & x"ff",
	4   => x"3018" & x"f0",
	5   => x"3034" & x"1a",
	6   => x"3035" & x"11",
	7   => x"3036" & x"69",
	8   => x"3037" & x"13",
	9   => x"3108" & x"01",
	10  => x"3630" & x"36",
	11  => x"3631" & x"0e",
	12  => x"3632" & x"e2",
	13  => x"3633" & x"12",
	14  => x"3621" & x"e0",
	15  => x"3704" & x"a0",
	16  => x"3703" & x"5a",
	17  => x"3715" & x"78",
	18  => x"3717" & x"01",
	19  => x"370b" & x"60",
	20  => x"3705" & x"1a",
	21  => x"3905" & x"02",
	22  => x"3906" & x"10",
	23  => x"3901" & x"0a",
	24  => x"3731" & x"12",
	25  => x"3600" & x"08",
	26  => x"3601" & x"33",
	27  => x"302d" & x"60",
	28  => x"3620" & x"52",
	29  => x"371b" & x"20",
	30  => x"471c" & x"50",
	31  => x"3a13" & x"43",
	32  => x"3a18" & x"00",
	33  => x"3a19" & x"f8",
	34  => x"3635" & x"13",
	35  => x"3636" & x"03",
	36  => x"3634" & x"40",
	37  => x"3622" & x"01",
	38  => x"3c01" & x"34",
	39  => x"3c04" & x"28",
	40  => x"3c05" & x"98",
	41  => x"3c06" & x"00",
	42  => x"3c07" & x"07",
	43  => x"3c08" & x"00",
	44  => x"3c09" & x"1c",
	45  => x"3c0a" & x"9c",
	46  => x"3c0b" & x"40",
	47  => x"3820" & x"42", 
	48  => x"3821" & x"02", 
	49  => x"3814" & x"11", 
	50  => x"3815" & x"11", 
	51  => x"3800" & x"01", 
	52  => x"3801" & x"50", 
	53  => x"3802" & x"01", 
	54  => x"3803" & x"b2", 
	55  => x"3804" & x"08", 
	56  => x"3805" & x"ef", 
	57  => x"3806" & x"05", 
	58  => x"3807" & x"f2", 
	59  => x"3808" & x"07", 
	60  => x"3809" & x"80", 
	61  => x"380a" & x"04", 
	62  => x"380b" & x"38", 
	63  => x"380c" & x"09", 
	64  => x"380d" & x"c4", 
	65  => x"380e" & x"04", 
	66  => x"380f" & x"60", 
	67  => x"3810" & x"00", 
	68  => x"3811" & x"10", 
	69  => x"3812" & x"00", 
	70  => x"3813" & x"04", 
	71  => x"3618" & x"04", 
	72  => x"3612" & x"2b", 
	73  => x"3708" & x"64", 
	74  => x"3709" & x"12", 
	75  => x"370c" & x"00", 
	76  => x"3a02" & x"04", 
	77  => x"3a03" & x"60", 
	78  => x"3a08" & x"01", 
	79  => x"3a09" & x"50", 
	80  => x"3a0a" & x"01", 
	81  => x"3a0b" & x"18", 
	82  => x"3a0e" & x"03", 
	83  => x"3a0d" & x"04", 
	84  => x"3a14" & x"04", 
	85  => x"3a15" & x"60", 
	86  => x"4001" & x"02", 
	87  => x"4004" & x"06", 
	88  => x"3000" & x"00", 
	89  => x"3001" & x"00", 
	90  => x"3002" & x"00", 
	91  => x"3004" & x"ff", 
	92  => x"3005" & x"ff", 
	93  => x"3006" & x"ff", 
	94  => x"3007" & x"ff", 
	95  => x"300e" & x"58", 
	96  => x"302e" & x"00", 
	97  => x"4740" & x"21", 
	98  => x"460b" & x"35", 
	99  => x"460c" & x"20", 
	100 => x"3824" & x"01", 
	101 => x"4300" & x"F8", 
	102 => x"5001" & x"01", 
	103 => x"501f" & x"03", 
	104 => x"5000" & x"06", 
	105 => x"5300" & x"08", 
	106 => x"5301" & x"30", 
	107 => x"5302" & x"10", 
	108 => x"5303" & x"00", 
	109 => x"5304" & x"08", 
	110 => x"5305" & x"30", 
	111 => x"5306" & x"08", 
	112 => x"5307" & x"16", 
	113 => x"5309" & x"08", 
	114 => x"530a" & x"30", 
	115 => x"530b" & x"04", 
	116 => x"530c" & x"06", 
	117 => x"5480" & x"01", 
	118 => x"5481" & x"08", 
	119 => x"5482" & x"14", 
	120 => x"5483" & x"28", 
	121 => x"5484" & x"51", 
	122 => x"5485" & x"65", 
	123 => x"5486" & x"71", 
	124 => x"5487" & x"7d", 
	125 => x"5488" & x"87", 
	126 => x"5489" & x"91", 
	127 => x"548a" & x"9a", 
	128 => x"548b" & x"aa", 
	129 => x"548c" & x"b8", 
	130 => x"548d" & x"cd", 
	131 => x"548e" & x"dd", 
	132 => x"548f" & x"ea", 
	133 => x"5490" & x"1d", 
	134 => x"5580" & x"02", 
	135 => x"5583" & x"40", 
	136 => x"5584" & x"10", 
	137 => x"5589" & x"10", 
	138 => x"558a" & x"00", 
	139 => x"558b" & x"f8", 
	140 => x"5800" & x"23", 
	141 => x"5801" & x"14", 
	142 => x"5802" & x"0f", 
	143 => x"5803" & x"0f", 
	144 => x"5804" & x"12", 
	145 => x"5805" & x"26", 
	146 => x"5806" & x"0c", 
	147 => x"5807" & x"08", 
	148 => x"5808" & x"05", 
	149 => x"5809" & x"05", 
	150 => x"580a" & x"08", 
	151 => x"580b" & x"0d", 
	152 => x"580c" & x"08", 
	153 => x"580d" & x"03", 
	154 => x"580e" & x"00", 
	155 => x"580f" & x"00", 
	156 => x"5810" & x"03", 
	157 => x"5811" & x"09", 
	158 => x"5812" & x"07", 
	159 => x"5813" & x"03", 
	160 => x"5814" & x"00", 
	161 => x"5815" & x"01", 
	162 => x"5816" & x"03", 
	163 => x"5817" & x"08", 
	164 => x"5818" & x"0d", 
	165 => x"5819" & x"08", 
	166 => x"581a" & x"05", 
	167 => x"581b" & x"06", 
	168 => x"581c" & x"08", 
	169 => x"581d" & x"0e", 
	170 => x"581e" & x"29", 
	171 => x"581f" & x"17", 
	172 => x"5820" & x"11", 
	173 => x"5821" & x"11", 
	174 => x"5822" & x"15", 
	175 => x"5823" & x"28", 
	176 => x"5824" & x"46", 
	177 => x"5825" & x"26", 
	178 => x"5826" & x"08", 
	179 => x"5827" & x"26", 
	180 => x"5828" & x"64", 
	181 => x"5829" & x"26", 
	182 => x"582a" & x"24", 
	183 => x"582b" & x"22", 
	184 => x"582c" & x"24", 
	185 => x"582d" & x"24", 
	186 => x"582e" & x"06", 
	187 => x"582f" & x"22", 
	188 => x"5830" & x"40", 
	189 => x"5831" & x"42", 
	190 => x"5832" & x"24", 
	191 => x"5833" & x"26", 
	192 => x"5834" & x"24", 
	193 => x"5835" & x"22", 
	194 => x"5836" & x"22", 
	195 => x"5837" & x"26", 
	196 => x"5838" & x"44", 
	197 => x"5839" & x"24", 
	198 => x"583a" & x"26", 
	199 => x"583b" & x"28", 
	200 => x"583c" & x"42", 
	201 => x"583d" & x"ce", 
	202 => x"5025" & x"00", 
	203 => x"3a0f" & x"30", 
	204 => x"3a10" & x"28", 
	205 => x"3a1b" & x"30", 
	206 => x"3a1e" & x"26", 
	207 => x"3a11" & x"60", 
	208 => x"3a1f" & x"14", 
	209 => x"4741" & x"00", 
	210 => x"3008" & x"02" 

	);

end ov5640_controller_pkg;