ibuf_inst : ibuf PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig
	);
